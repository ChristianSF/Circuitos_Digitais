module porta_not_verilog (a, b);
input wire a;
output wire b;

assign b = ~a;

endmodule
