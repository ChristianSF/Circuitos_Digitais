module exemplo_AND(A, B, C);
input wire A, B;
output wire C;

assign C = A & B;

endmodule
